module Buzzer2 (
    input wire clk,         // Clock signal
    input wire [3:0] note,
    input enable,
    output wire speaker     // Buzzer output signal
) ;

    wire [31:0] notes [7:0];
    reg [31:0] counter;
    reg pwm;

    // Frequencies of do , re , mi , fa , so , la , si
    // Obtain the ratio of how long the buzzer should be active in one second
    assign notes[1] = 381680;
    assign notes[2] = 340136;
    assign notes[3] = 303030;
    assign notes[4] = 285714;
    assign notes[5] = 255102;
    assign notes[6] = 227273;
    assign notes[7] = 202429;
    
    initial begin
        pwm = 0;
    end

    always @ ( posedge clk ) begin
        if(enable==1'b0)
            pwm<=0;
        else if (counter < notes [note] || note == 1'b0) begin
            counter <= counter + 1'b1;
        end 
        else begin
            pwm = ~pwm;
            counter <= 0;
        end
    end

    assign speaker = pwm; // Output a PWM signal to the buzzer
    
endmodule